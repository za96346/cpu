module Top_pipeline(
    input logic clk;
    input logic reset;
);
    
endmodule